-----------------------------
--PROGETTO FFT 16x16
--AMATO GIOVANNI LUCA Matr.267511
--CERBAI MATILDE Matr.274908 
--CHISCIOTTI LAURA Matr.274728
--GOTI GIANLUCA Matr.269825
-----------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mux3dp is
	generic ( parallelism: integer := 24 );
port(
	d1: in signed(parallelism-1 downto 0);
	d2: in signed(parallelism*2 downto 0);
	q: out signed(parallelism*2 downto 0);
	sel: in std_logic
	);
end mux3dp;

architecture behavioural of mux3dp is
		begin
			mux_proc:process(d1,d2,sel)
			begin
				case sel is
					when '0' =>
						
						q<=shift_left(resize(d1,49),25); 

					when others =>
						q<=d2;
				end case;
			end process mux_proc;
	end behavioural;
			